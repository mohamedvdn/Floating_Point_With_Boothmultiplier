module Main_Adder_Tree(PP0,PP1,PP2,PP3,PP4,PP5,PP6,PP7,P);
  input [63:0]PP0;
  input [63:0]PP1; 
  input [63:0]PP2;  
  input [63:0]PP3;  
  input [63:0]PP4;    
  input [63:0]PP5;    
  input [63:0]PP6;    
  input [63:0]PP7;    
  
  output [63:0]P;
  
  wire [4:0]W4,W5,W6,W7,W8,W9,W10,W11,W12,W13,W14,W15,W16,W17,W18,W19,W20,W21,W22,W23,W24,W25,W26,W27,W28,W29,W30,W31,W32,W33,W34,W35,W36,W37,W38,W39,W40,W41,W42,W43,W44,W45,W46,W47,W48,W49,W50,W51,W52,W53,W54,W55,W56,W57,W58,W59,W60,W61,W62;
  
       assign P[0]=PP0[0];
       assign P[1]=PP0[1];
       assign P[2]=PP0[2];
       assign P[3]=PP0[3];  
  assign {W4,P[4]}=PP0[4]+PP1[0];
  assign {W5,P[5]}=PP0[5]+PP1[1]+W4;
  assign {W6,P[6]}=PP0[6]+PP1[2]+W5;
  assign {W7,P[7]}=PP0[7]+PP1[3]+W6;        
  assign {W8,P[8]}=PP0[8]+PP1[4]+PP2[0]+W7;        
  assign {W9,P[9]}=PP0[9]+PP1[5]+PP2[1]+W8;        
assign {W10,P[10]}=PP0[10]+PP1[6]+PP2[2]+W9;        
assign {W11,P[11]}=PP0[11]+PP1[7]+PP2[3]+W10;        
assign {W12,P[12]}=PP0[12]+PP1[8]+PP2[4]+PP3[0]+W11;        
assign {W13,P[13]}=PP0[13]+PP1[9]+PP2[5]+PP3[1]+W12;         
assign {W14,P[14]}=PP0[14]+PP1[10]+PP2[6]+PP3[2]+W13;         
assign {W15,P[15]}=PP0[15]+PP1[11]+PP2[7]+PP3[3]+W14;         
assign {W16,P[16]}=PP0[16]+PP1[12]+PP2[8]+PP3[4]+PP4[0]+W15;         
assign {W17,P[17]}=PP0[17]+PP1[13]+PP2[9]+PP3[5]+PP4[1]+W16;         
assign {W18,P[18]}=PP0[18]+PP1[14]+PP2[10]+PP3[6]+PP4[2]+W17;           
assign {W19,P[19]}=PP0[19]+PP1[15]+PP2[11]+PP3[7]+PP4[3]+W18;           
assign {W20,P[20]}=PP0[20]+PP1[16]+PP2[12]+PP3[8]+PP4[4]+PP5[0]+W19;             
assign {W21,P[21]}=PP0[21]+PP1[17]+PP2[13]+PP3[9]+PP4[5]+PP5[1]+W20;             
assign {W22,P[22]}=PP0[22]+PP1[18]+PP2[14]+PP3[10]+PP4[6]+PP5[2]+W21;               
assign {W23,P[23]}=PP0[23]+PP1[19]+PP2[15]+PP3[11]+PP4[7]+PP5[3]+W22;               
assign {W24,P[24]}=PP0[24]+PP1[20]+PP2[16]+PP3[12]+PP4[8]+PP5[4]+PP6[0]+W23;               
assign {W25,P[25]}=PP0[25]+PP1[21]+PP2[17]+PP3[13]+PP4[9]+PP5[5]+PP6[1]+W24;                 
assign {W26,P[26]}=PP0[26]+PP1[22]+PP2[18]+PP3[14]+PP4[10]+PP5[6]+PP6[2]+W25;                 
assign {W27,P[27]}=PP0[27]+PP1[23]+PP2[19]+PP3[15]+PP4[11]+PP5[7]+PP6[3]+W26;                   
assign {W28,P[28]}=PP0[28]+PP1[24]+PP2[20]+PP3[16]+PP4[12]+PP5[8]+PP6[4]+PP7[0]+W27;                   
assign {W29,P[29]}=PP0[29]+PP1[25]+PP2[21]+PP3[17]+PP4[13]+PP5[9]+PP6[5]+PP7[1]+W28;                   
assign {W30,P[30]}=PP0[30]+PP1[26]+PP2[22]+PP3[18]+PP4[14]+PP5[10]+PP6[6]+PP7[2]+W29;                   
assign {W31,P[31]}=PP0[31]+PP1[27]+PP2[23]+PP3[19]+PP4[15]+PP5[11]+PP6[7]+PP7[3]+W30;                   
assign {W32,P[32]}=PP0[32]+PP1[28]+PP2[24]+PP3[20]+PP4[16]+PP5[12]+PP6[8]+PP7[4]+W31;                   
assign {W33,P[33]}=PP0[33]+PP1[29]+PP2[25]+PP3[21]+PP4[17]+PP5[13]+PP6[9]+PP7[5]+W32;                   
assign {W34,P[34]}=PP0[34]+PP1[30]+PP2[26]+PP3[22]+PP4[18]+PP5[14]+PP6[10]+PP7[6]+W33;                   
assign {W35,P[35]}=PP0[35]+PP1[31]+PP2[27]+PP3[23]+PP4[19]+PP5[15]+PP6[11]+PP7[7]+W34;                   
assign {W36,P[36]}=PP0[36]+PP1[32]+PP2[28]+PP3[24]+PP4[20]+PP5[16]+PP6[12]+PP7[8]+W35;                   
assign {W37,P[37]}=PP0[37]+PP1[33]+PP2[29]+PP3[25]+PP4[21]+PP5[17]+PP6[13]+PP7[9]+W36;                   
assign {W38,P[38]}=PP0[38]+PP1[34]+PP2[30]+PP3[26]+PP4[22]+PP5[18]+PP6[14]+PP7[10]+W37;                   
assign {W39,P[39]}=PP0[39]+PP1[35]+PP2[31]+PP3[27]+PP4[23]+PP5[19]+PP6[15]+PP7[11]+W38;                   
assign {W40,P[40]}=PP0[40]+PP1[36]+PP2[32]+PP3[28]+PP4[24]+PP5[20]+PP6[16]+PP7[12]+W39;                   
assign {W41,P[41]}=PP0[41]+PP1[37]+PP2[33]+PP3[29]+PP4[25]+PP5[21]+PP6[17]+PP7[13]+W40;                   
assign {W42,P[42]}=PP0[42]+PP1[38]+PP2[34]+PP3[30]+PP4[26]+PP5[22]+PP6[18]+PP7[14]+W41;                   
assign {W43,P[43]}=PP0[43]+PP1[39]+PP2[35]+PP3[31]+PP4[27]+PP5[23]+PP6[19]+PP7[15]+W42;                   
assign {W44,P[44]}=PP0[44]+PP1[40]+PP2[36]+PP3[32]+PP4[28]+PP5[24]+PP6[20]+PP7[16]+W43;                   
assign {W45,P[45]}=PP0[45]+PP1[41]+PP2[37]+PP3[33]+PP4[29]+PP5[25]+PP6[21]+PP7[17]+W44;                   
assign {W46,P[46]}=PP0[46]+PP1[42]+PP2[38]+PP3[34]+PP4[30]+PP5[26]+PP6[22]+PP7[18]+W45;                   
assign {W47,P[47]}=PP0[47]+PP1[43]+PP2[39]+PP3[35]+PP4[31]+PP5[27]+PP6[23]+PP7[19]+W46;                   
assign {W48,P[48]}=PP0[48]+PP1[44]+PP2[40]+PP3[36]+PP4[32]+PP5[28]+PP6[24]+PP7[20]+W47;                   
assign {W49,P[49]}=PP0[49]+PP1[45]+PP2[41]+PP3[37]+PP4[33]+PP5[29]+PP6[25]+PP7[21]+W48;                   
assign {W50,P[50]}=PP0[50]+PP1[46]+PP2[42]+PP3[38]+PP4[34]+PP5[30]+PP6[26]+PP7[22]+W49;                   
assign {W51,P[51]}=PP0[51]+PP1[47]+PP2[43]+PP3[39]+PP4[35]+PP5[31]+PP6[27]+PP7[23]+W50;                   
assign {W52,P[52]}=PP0[52]+PP1[48]+PP2[44]+PP3[40]+PP4[36]+PP5[32]+PP6[28]+PP7[24]+W51;                   
assign {W53,P[53]}=PP0[53]+PP1[49]+PP2[45]+PP3[41]+PP4[37]+PP5[33]+PP6[29]+PP7[25]+W52;                   
assign {W54,P[54]}=PP0[54]+PP1[50]+PP2[46]+PP3[42]+PP4[38]+PP5[34]+PP6[30]+PP7[26]+W53;                   
assign {W55,P[55]}=PP0[55]+PP1[51]+PP2[47]+PP3[43]+PP4[39]+PP5[35]+PP6[31]+PP7[27]+W54;                   
assign {W56,P[56]}=PP0[56]+PP1[52]+PP2[48]+PP3[44]+PP4[40]+PP5[36]+PP6[32]+PP7[28]+W55;                   
assign {W57,P[57]}=PP0[57]+PP1[53]+PP2[49]+PP3[45]+PP4[41]+PP5[37]+PP6[33]+PP7[29]+W56;                   
assign {W58,P[58]}=PP0[58]+PP1[54]+PP2[50]+PP3[46]+PP4[42]+PP5[38]+PP6[34]+PP7[30]+W57;                   
assign {W59,P[59]}=PP0[59]+PP1[55]+PP2[51]+PP3[47]+PP4[43]+PP5[39]+PP6[35]+PP7[31]+W58;                   
assign {W60,P[60]}=PP0[60]+PP1[56]+PP2[52]+PP3[48]+PP4[44]+PP5[40]+PP6[36]+PP7[32]+W59;                   
assign {W61,P[61]}=PP0[61]+PP1[57]+PP2[53]+PP3[49]+PP4[45]+PP5[41]+PP6[37]+PP7[33]+W60;                   
assign {W62,P[62]}=PP0[62]+PP1[58]+PP2[54]+PP3[50]+PP4[46]+PP5[42]+PP6[38]+PP7[34]+W61;                   
assign {W63,P[63]}=PP0[63]+PP1[59]+PP2[55]+PP3[51]+PP4[47]+PP5[43]+PP6[39]+PP7[35]+W62;                   


endmodule