module M_white_ball (A,B,C,D);
input A,B;  
output C,D; 
and m1 (C,A,A);
and m2 (D,B,B);
endmodule 