library verilog;
use verilog.vl_types.all;
entity Floating_Point_Multiplier_Vedic_hybrid_Tb is
end Floating_Point_Multiplier_Vedic_hybrid_Tb;
